//Compuerta AND

module Compuerta_and(
	input [3:0] A,
	input [3:0] B,
	output [3:0] F
	);

assign F = A & B;
endmodule
