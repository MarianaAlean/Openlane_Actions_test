//Compuerta NOT

module Compuerta_not(
	input [3:0] A,
	output [3:0] F
	);

assign F = ~A;
endmodule
