//Comparador >

module mayor(
	input [3:0] A,
	input [3:0] B,
	output F
	);

assign F = (A > B);

endmodule
